/Users/gunwoo/.dotfiles/vim/bundle/ale/test/test-files/hdl_server/with_config_file/foo.vhd