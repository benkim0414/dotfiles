/Users/gunwoo/.dotfiles/vim/bundle/ale/test/test-files/hdl_server/with_git/files/foo.vhd