/Users/gunwoo/.dotfiles/vim/bundle/ale/test/test-files/hdl_server/foo.vhd